`timescale 1ns / 1ps

module main(
  input sys_clk,
  input rst_n,
);

endmodule
