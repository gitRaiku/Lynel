`timescale 1ns / 1ps

`include usb.v


module ();

endmodule
