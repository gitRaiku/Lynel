module usb(

);

endmodule
