../usbi2c.srcs/sources_1/new/cdc.sv